module enet(ENET_DATA, ENET_CLK, ENET_CMD, ENET_CS_N, ENET_INT, ENET_RD_N, ENET_WR_N, ENET_RST_N);
	input [15:0] ENET_DATA;
	input ENET_CLK;
	input ENET_CMD;
	input ENET_CS_N;
	input ENET_INT;
	input ENET_RD_N;
	input ENET_WR_N;
	input ENET_RST_N;
endmodule 